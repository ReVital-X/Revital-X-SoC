`timescale 1ns / 1ps
module instruction_fetch(
    input clk,rst,
    output reg [31:0]pc
    );
    
    always @(posedge clk or posedge rst) begin
        if(rst)
            pc <= 32'h0;
            
        else
            pc <= pc + 4;
    end
    
endmodule
